interface calculator_inter;

  logic [7:0] a;
  logic [7:0] b;
  logic [7:0] result;
  logic [2:0] opcode;

endinterface

